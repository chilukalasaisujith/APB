`ifndef _con_
`define _con_

class configuration;
int txn_num;
endclass
`endif
`ifndef  base
`define  base

class base;
rand bit [3:0]addr;
rand bit [7:0]data;
bit write;
bit [7:0]read_data;
bit [7:0] exp_read_data;
endclass

`endif